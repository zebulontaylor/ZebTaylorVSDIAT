magic
tech sky130A
magscale 1 2
timestamp 1753113566
<< error_p >>
rect 2706 2412 2720 2414
rect 1260 1970 1274 2220
rect 1920 2052 1940 2342
rect 2748 1970 2762 2412
rect 3198 2032 3226 2444
rect 3464 2038 3502 2464
rect 3754 2050 3792 2476
rect 4226 2462 4233 2598
rect 5003 2570 5006 2581
rect 5014 2474 5021 2570
rect 4224 2154 4233 2314
rect 5001 2254 5006 2265
rect 5012 2158 5021 2254
rect 1780 978 1790 1292
rect 3012 1288 3058 1302
rect 2508 962 2534 1276
rect 3638 896 3640 1308
rect 4949 940 4950 941
rect 4950 939 4951 940
rect 5538 926 5539 927
rect 5537 925 5538 926
rect 5530 894 5531 895
rect 5529 893 5530 894
rect 3004 738 3050 752
rect 1768 398 1778 712
rect 2496 382 2522 696
rect 5560 506 5561 507
rect 5559 505 5560 506
rect 5552 474 5553 475
rect 5551 473 5552 474
rect 4917 434 4918 435
rect 4918 433 4919 434
rect 2718 22 2980 104
rect 3062 22 3326 98
rect 2606 -426 2608 -14
rect 3988 -16 4222 46
rect 4238 -16 4500 68
rect 4582 -16 4804 62
rect 2814 -420 2884 -364
rect 3158 -426 3230 -364
rect 4126 -462 4128 -50
rect 4334 -456 4404 -400
rect 4678 -462 4750 -400
<< nwell >>
rect 1554 2556 2344 2558
rect 1554 1794 2462 2556
rect 4042 2410 5440 2752
rect 2178 1792 2462 1794
rect 1586 824 3232 1414
rect 4566 1150 5554 1152
rect 4566 720 5780 1150
rect 5202 718 5780 720
rect 3848 -90 4880 146
rect 3930 -694 4874 -346
<< nmos >>
rect 1732 398 1778 712
rect 2546 382 2592 696
rect 3004 412 3050 726
rect 5560 506 5592 558
rect 4830 434 4918 486
rect 4830 352 4962 434
rect 5520 474 5592 506
rect 5520 416 5552 474
<< pmos >>
rect 1744 978 1790 1292
rect 2558 962 2604 1276
rect 3012 962 3058 1276
rect 4862 940 4950 992
rect 4862 858 4994 940
rect 5538 926 5570 978
rect 5498 894 5570 926
rect 5498 836 5530 894
<< pmoslvt >>
rect 1870 2052 1920 2342
<< ndiff >>
rect 4224 2154 4434 2314
rect 1670 398 1732 712
rect 1778 398 1828 712
rect 2522 382 2546 696
rect 2592 382 2644 696
rect 2952 412 3004 726
rect 3050 412 3102 726
rect 5468 506 5560 558
rect 4778 352 4830 486
rect 4962 352 5014 434
rect 5468 416 5520 506
rect 5592 474 5704 558
rect 5552 416 5704 474
rect 2498 -590 3310 -460
<< pdiff >>
rect 1730 2052 1870 2342
rect 1920 2052 2012 2342
rect 4226 2462 4438 2598
rect 1682 978 1744 1292
rect 1790 978 1840 1292
rect 2534 962 2558 1276
rect 2604 962 2656 1276
rect 2960 962 3012 1276
rect 3058 962 3110 1276
rect 4810 858 4862 992
rect 4994 858 5046 940
rect 5446 926 5538 978
rect 5446 836 5498 926
rect 5570 894 5682 978
rect 5530 836 5682 894
rect 4016 -626 4828 -496
<< psubdiff >>
rect 5012 2158 5182 2254
rect 1828 604 2166 712
rect 1828 492 2036 604
rect 2144 492 2166 604
rect 1828 398 2166 492
rect 4600 482 4664 506
rect 4600 394 4664 418
rect 5236 480 5300 504
rect 5236 392 5300 416
rect 2534 22 3350 118
<< nsubdiff >>
rect 2248 2230 2408 2270
rect 2248 2040 2408 2076
rect 4640 2540 4704 2564
rect 4640 2452 4704 2476
rect 5014 2474 5184 2570
rect 1840 1184 2178 1292
rect 1840 1072 2048 1184
rect 2156 1072 2178 1184
rect 1840 978 2178 1072
rect 4632 988 4696 1012
rect 4632 900 4696 924
rect 5268 986 5332 1010
rect 5268 898 5332 922
rect 3988 -16 4804 80
<< psubdiffcont >>
rect 2036 492 2144 604
rect 4600 418 4664 482
rect 5236 416 5300 480
<< nsubdiffcont >>
rect 2248 2076 2408 2230
rect 4640 2476 4704 2540
rect 2048 1072 2156 1184
rect 4632 924 4696 988
rect 5268 922 5332 986
<< poly >>
rect 1870 2342 1920 2452
rect 1244 1970 1260 2220
rect 1870 1946 1920 2052
rect 2638 1970 2720 2414
rect 2748 1968 2830 2412
rect 4140 2062 4218 2759
rect 4928 2076 5006 2789
rect 1744 1292 1790 1360
rect 2558 1276 2604 1344
rect 3012 1276 3058 1288
rect 1744 928 1790 978
rect 2558 912 2604 962
rect 3012 912 3058 962
rect 4862 992 4994 1018
rect 4950 940 4994 992
rect 5538 978 5570 1016
rect 1732 712 1778 780
rect 2546 696 2592 764
rect 3004 726 3050 738
rect 1732 348 1778 398
rect 3544 708 4304 854
rect 4862 808 4994 858
rect 5498 806 5530 836
rect 5560 558 5592 596
rect 4830 486 4962 512
rect 2546 332 2592 382
rect 3004 362 3050 412
rect 4918 434 4962 486
rect 5520 386 5552 416
rect 4830 302 4962 352
<< npolyres >>
rect 3160 2032 3198 2444
rect 3574 896 3638 1308
rect 2542 -426 2606 -14
rect 4062 -462 4126 -50
<< ppolyres >>
rect 3432 2038 3464 2464
rect 3846 902 3916 1330
rect 2814 -420 2884 8
rect 4334 -456 4404 -28
<< xpolyres >>
rect 3722 2050 3754 2476
rect 4190 896 4262 1324
rect 3158 -426 3230 2
rect 4678 -462 4750 -34
<< locali >>
rect 4640 2540 4704 2564
rect 4640 2452 4704 2476
rect 2248 2230 2408 2270
rect 2248 2040 2408 2076
rect 2048 1184 2156 1204
rect 2048 1046 2156 1072
rect 4632 988 4696 1012
rect 4632 900 4696 924
rect 5268 986 5332 1010
rect 5268 898 5332 922
rect 2036 604 2144 624
rect 2036 466 2144 492
rect 4600 482 4664 506
rect 4600 394 4664 418
rect 5236 480 5300 504
rect 5236 392 5300 416
<< labels >>
flabel comment s 292 2248 292 2248 0 FreeSans 800 0 0 0 Poly
flabel comment s 1878 1862 1878 1862 0 FreeSans 560 0 0 0 poly.1b
flabel comment s 1272 1850 1272 1850 0 FreeSans 560 0 0 0 poly.1a
flabel comment s 2766 1836 2766 1842 0 FreeSans 560 0 0 0 poly.2
flabel comment s 3482 1892 3482 1894 0 FreeSans 560 0 0 0 poly.3
flabel comment s 4264 1904 4264 1904 0 FreeSans 560 0 0 0 poly.4
flabel comment s 5030 1944 5030 1944 0 FreeSans 560 0 0 0 poly.5
flabel comment s 5088 2338 5088 2338 0 FreeSans 560 0 0 0 Incorrect_flags_poly.4
flabel comment s 484 1360 490 1360 0 FreeSans 560 0 0 0 Correct_by_design
flabel comment s 1874 236 1874 242 0 FreeSans 560 0 0 0 poly.6
flabel comment s 2612 244 2612 250 0 FreeSans 560 0 0 0 poly.7
flabel comment s 3090 248 3090 254 0 FreeSans 560 0 0 0 poly.8
flabel comment s 3916 482 3916 488 0 FreeSans 560 0 0 0 poly.9
flabel comment s 3886 610 3886 610 0 FreeSans 560 0 0 0 Incorrect
flabel comment s 4792 200 4792 200 0 FreeSans 560 0 0 0 poly.10
flabel comment s 5428 198 5428 198 0 FreeSans 560 0 0 0 poly.11
flabel comment s 410 1196 410 1196 0 FreeSans 560 0 0 0 poly.12
flabel comment s 376 1026 376 1026 0 FreeSans 560 0 0 0 poly.15
flabel comment s 408 552 408 552 0 FreeSans 560 0 0 0 Not implemented
flabel comment s 476 334 476 334 0 FreeSans 560 0 0 0 poly.16
<< end >>
