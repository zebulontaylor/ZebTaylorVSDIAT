magic
tech sky130A
magscale 1 2
timestamp 1753112212
<< error_p >>
rect 2679 2239 2688 2248
rect 2670 2230 2673 2239
rect 2670 2183 2673 2192
rect 2679 2174 2688 2183
rect 3243 980 3264 1435
rect 3303 1040 3344 1375
<< metal2 >>
rect 2673 2183 2679 2239
rect 2739 2183 2795 2239
<< via2 >>
rect 2679 2183 2739 2239
<< metal3 >>
rect 1418 2250 1716 2328
rect 1419 2248 1715 2250
rect 2092 2140 2432 2302
rect 2679 2266 2739 2376
rect 2674 2248 2744 2266
rect 2666 2239 2748 2248
rect 2666 2183 2679 2239
rect 2739 2183 2748 2239
rect 2666 2174 2748 2183
rect 3068 2174 3190 2286
rect 1449 1461 2149 1583
rect 1375 1398 2149 1461
rect 1449 1338 2149 1398
rect 1375 1275 2149 1338
rect 1449 883 2149 1275
rect 2564 866 3264 1566
rect 3303 1040 3380 1375
<< labels >>
flabel comment s 1791 1664 1791 1664 0 FreeSans 560 0 0 0 Not implemented
flabel comment s 1549 2081 1549 2081 0 FreeSans 560 0 0 0 m3.1
flabel comment s 2260 2050 2260 2050 0 FreeSans 560 0 0 0 m3.2
flabel comment s 2974 811 2974 811 0 FreeSans 560 0 0 0 m3.3d
flabel comment s 1821 811 1821 811 0 FreeSans 560 0 0 0 m3.3c
flabel comment s 2712 2108 2712 2108 0 FreeSans 560 0 0 0 m3.5
flabel comment s 3131 2080 3131 2080 0 FreeSans 560 0 0 0 m3.6
flabel comment s 700 2120 700 2120 0 FreeSans 560 0 0 0 Correct by design
flabel comment s 688 2342 688 2342 0 FreeSans 800 0 0 0 Met3 (m3)
flabel comment s 725 1999 725 1999 0 FreeSans 560 0 0 0 m3.4
<< end >>
